magic
tech sky130A
magscale 1 2
timestamp 1741220675
<< checkpaint >>
rect -1549 6296 2491 6304
rect -1549 5960 2492 6296
rect -1549 5540 2760 5960
rect -1664 -2186 2992 5540
<< error_s >>
rect 160 2132 166 2138
rect 154 2126 160 2132
rect 154 2068 160 2074
rect 160 2062 166 2068
<< locali >>
rect -200 710 -8 954
rect 952 710 1144 996
rect -300 690 1206 710
rect -300 510 190 690
rect 370 510 1206 690
rect -300 500 1206 510
<< viali >>
rect 190 510 370 690
<< metal1 >>
rect -1 4599 0 4601
rect 200 4500 300 4689
rect 700 4600 1000 4700
rect 700 4500 800 4600
rect 62 3038 115 4500
rect 56 3032 120 3038
rect 50 2968 56 3032
rect 120 2968 126 3032
rect 56 2962 120 2968
rect 62 974 115 2962
rect 184 690 376 4500
rect 900 3900 1000 4600
rect 1299 4499 1301 4500
rect 700 3800 1000 3900
rect 700 3700 800 3800
rect 668 3032 732 3038
rect 662 2968 668 3032
rect 732 2968 738 3032
rect 668 2962 732 2968
rect 900 2300 1000 3800
rect 700 2200 1000 2300
rect 700 2100 800 2200
rect 900 1500 1000 2200
rect 700 1400 1000 1500
rect 700 1300 800 1400
rect 900 800 1000 1400
rect 184 510 190 690
rect 370 510 376 690
rect 184 498 376 510
<< via1 >>
rect 56 2968 120 3032
rect 668 2968 732 3032
<< metal2 >>
rect 56 3032 120 3038
rect 50 2968 56 3032
rect 56 2932 120 2968
rect 668 3032 732 3038
rect 732 2968 738 3032
rect 668 2932 732 2968
rect 56 2868 732 2932
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 -104 0 1 4001
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1740610800
transform 1 0 -104 0 1 802
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1740610800
transform 1 0 -104 0 1 1601
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1740610800
transform 1 0 -104 0 1 2403
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_4
timestamp 1740610800
transform 1 0 -104 0 1 3200
box -184 -128 1336 928
<< labels >>
flabel metal1 700 4500 800 4700 0 FreeSans 1600 0 0 0 IBNS_20U
port 1 nsew
flabel locali -300 500 190 710 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel metal2 56 2868 732 2932 0 FreeSans 1600 0 0 0 IBPS_5U
port 5 nsew
<< end >>
